interface muxi;
  logic a,b,c,d,e,f,g,h;
  logic [2:0]sel;
  logic yout;
endinterface
