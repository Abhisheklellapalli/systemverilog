module subtraction(input [2:0]a,b,output [2:0]sub);
  assign sub = a-b;
endmodule
