interface fa;
  logic a,b;
  logic sum,cout;
endinterface
